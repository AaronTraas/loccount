//Hello, World in Verilog
module top;

initial
    $display("Hello, world!");

endmodule
